* EESchema Netlist Version 1.1 (Spice format) creation date: 6/4/2009-01:47:07


U4  N-000017 N-000002 N-000014 VCC PHDARL
U3  N-000005 N-000019 GND N-000009 PHDARL
U2  N-000006 N-000002 N-000010 VCC PHDARL
U1  N-000016 N-000018 GND N-000015 PHDARL
P3  N-000013 N-000004 CONN_2
P2  GND VCC CONN_2
Q4  GND N-000011 N-000013 NPN
Q2  GND N-000007 N-000004 NPN
Q3  VCC N-000012 N-000013 PNP
Q1  VCC N-000008 N-000004 PNP
K1  N-000002 N-000018 N-000019 CONN_3
R9  VCC N-000008 10k
R11  VCC N-000012 10k
R10  N-000007 GND 10k
R12  N-000011 GND 10k
R8  N-000014 N-000011 1k
R7  N-000009 N-000012 1k
R5  N-000008 N-000015 1k
R6  N-000007 N-000010 1k
R1  N-000016 N-000019 470
R2  N-000006 N-000018 470
R4  N-000019 N-000017 470
R3  N-000018 N-000005 470

.end
